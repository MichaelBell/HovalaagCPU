`timescale 1ns / 1ps
// Copyright (C) 2020 Michael Bell

// Insert the program output by the 'bintoverilog.py' script below.
module Program(
    input clk,
    input [7:0] addr,
    output reg [31:0] data
    );

		//8'h00:   data = 32'b00000011000000000000000001000000;
		//8'h01:   data = 32'b01010100000010001100000000000001;

	always @(posedge clk) begin
		case (addr)     //  ALU-A-B-C-DW-F-PCOIXK-----L-----
		8'h00:   data = 32'b00000011000000100001000010011111;
		8'h01:   data = 32'b00100011010000000001000000001010;
		8'h02:   data = 32'b00100111000000000001000000001111;
		8'h03:   data = 32'b00100111001000001000010001000100;
		8'h04:   data = 32'b00000000000010000001000000000000;
		8'h05:   data = 32'b00010000000010000101000000000000;
		8'h06:   data = 32'b00100000000010000101000000000000;
		8'h07:   data = 32'b00110000000010000101000000000000;
		8'h08:   data = 32'b01000000000010000101000000000000;
		8'h09:   data = 32'b01010000000010000101000000000000;
		8'h0a:   data = 32'b01100000000010000101000000000000;
		8'h0b:   data = 32'b01110000000010000101000000000000;
		8'h0c:   data = 32'b10000000000010000101000000000000;
		8'h0d:   data = 32'b10100000000010000101000000000000;
		8'h0e:   data = 32'b10010000000010000101000000000000;
		8'h0f:   data = 32'b10110000000010000101000000000000;
		8'h10:   data = 32'b11000000000010000101000000000000;
		8'h11:   data = 32'b00001000001000001101000000000100;


		
		default: data = 32'b00000000000000001000000000000000;
		endcase
	end

endmodule
